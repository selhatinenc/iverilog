module helloword;
	initial begin
		$display("Hello word!");
	end
endmodule;