module  test(
    
);

    
endmodule