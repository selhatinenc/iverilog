module dff_sync_res(D, clk, sync_reset, Q);
    input D;
    input clk;
    input sync_reset;
    output reg Q;

    always @(posedge clk)
    begin
        if(sync_reset==1)
            Q <= 0;
        else    
            Q<=D;
    end

    // Your code goes here.  DO NOT change anything that is already given! Otherwise, you will not be able to pass the tests!

endmodule 